system_pll_inst : system_pll PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
